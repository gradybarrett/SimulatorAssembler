"0011000000001001"  -- 0: store a 9
"0011010000001010"  -- 1: store b 10
"0101100000001001"  -- 2: seti c 9
"0101110000001010"  -- 3: seti d 10
"1000001000000000"  -- 4: addptr a c 0
"1000001100000000"  -- 5: addptr a d 0
"1000001000000001"  -- 6: addptr a c 1
"1011001000000000"  -- 7: storeptr a c 0
"1011001100000000"  -- 8: storeptr a d 0
"1011001000000001"  -- 9: storeptr a c 1
"1001001000000000"  -- 10: subptr a c 0
"1001001100000000"  -- 11: subptr a d 0
"1001001000000001"  -- 12: subptr a c 1
"1010001000000000"  -- 13: loadptr a c 0
"1010001100000000"  -- 14: loadptr a d 0
"1010001000000001"  -- 15: loadptr a c 1
