"0100000000000001"  -- 0: addi a 1
"0000010000000001"  -- 1: add b 1
"1000100000000000"  -- 2: addptr c a 0
"1000110000000010"  -- 3: addptr d a 2
"0101000000000000"  -- 4: seti a 0
"0001010000000001"  -- 5: sub b 1
"0101000000000011"  -- 6: seti a 3
"0101010000000100"  -- 7: seti b 4
"1001010000000000"  -- 8: subptr b a 0
"0111000000001000"  -- 9: jz a 8
"0110000000000001"  -- 10: jump 1
"0101000000000000"  -- 11: seti a 0
"1010010000000000"  -- 12: loadptr b a 0
"0100000000001010"  -- 13: addi a 10
"1011000100000000"  -- 14: storeptr a b 0
