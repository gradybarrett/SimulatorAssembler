"0101000000000011"  -- 0: seti a 3
"0111000000000101"  -- 1: jz a 5
"0001000000000010"  -- 2: sub a 2
"0100000000000001"  -- 3: addi a 1
"0110000000000001"  -- 4: jump 1
"0011000000000000"  -- 6: store a 0
"0011000000001001"  -- 7: store a 9
"0011010000001010"  -- 8: store b 10
"0101000000000000"  -- 9: seti a 0
"0101010000000000"  -- 10: seti b 0
"0001010000000001"  -- 11: sub b 1
"0101100000001001"  -- 12: seti c 9
"0101110000001010"  -- 13: seti d 10
"1000000000000000"  -- 14: addptr a a 0
"1000000100000000"  -- 15: addptr a b 0
"1000001000000000"  -- 16: addptr a c 0
"1000001100000000"  -- 17: addptr a d 0
"1000001000000001"  -- 18: addptr a c 1
"1011000000000000"  -- 19: storeptr a a 0
"1011000100000000"  -- 20: storeptr a b 0
"1011001000000000"  -- 21: storeptr a c 0
"1011001100000000"  -- 22: storeptr a d 0
"1011001000000001"  -- 23: storeptr a c 1
"1001000000000000"  -- 24: subptr a a 0
"1001000100000000"  -- 25: subptr a b 0
"1001001000000000"  -- 26: subptr a c 0
"1001001100000000"  -- 27: subptr a d 0
"1001001000000001"  -- 28: subptr a c 1
"1010000000000000"  -- 29: loadptr a a 0
"1010000100000000"  -- 30: loadptr a b 0
"1010001000000000"  -- 31: loadptr a c 0
"1010001100000000"  -- 32: loadptr a d 0
"1010001000000001"  -- 33: loadptr a c 1
"0010000000000000"  -- 34: load a 0
"0010010000000101"  -- 35: load b 5
"0010100000001001"  -- 36: load c 9
"0010110000001010"  -- 37: load d 10
"0000000000000000"  -- 39: add a 0
"0000010000001001"  -- 40: add b 9
"0000010000001010"  -- 41: add b 10
"0001000000000000"  -- 42: sub a 0
"0001010000001001"  -- 43: sub b 9
"0001010000001010"  -- 44: sub b 10
"0110000000101011"  -- 45: jump 43
"0101100001100011"  -- 46: seti c 99
"0101110001100011"  -- 47: seti d 99
